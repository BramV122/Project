module Project();


endmodule 